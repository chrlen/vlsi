-- Schnittstelle der Testbench

library IEEE;
use IEEE.std_logic_1164.all;

LIBRARY work;
use work.delayPack.ALL;

ENTITY func_tb IS
END func_tb;
