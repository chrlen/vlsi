configuration dummy_mhdl_cfg_FUNC_TB of FUNC_TB is
for ARCH
end for;
end;
